module slave (
    input CS,   // chip select from master
    input SCLK, // SPI clock (the driven one)
    input SDI,  // slave data in (from master)
    //
    output SDO  // slave data out (to master)
);



endmodule