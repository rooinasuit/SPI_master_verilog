interface m_int();

logic [7:0] MOSI_data;
logic MISO;
logic [7:0] MISO_data;
logic [7:0] master_stash_ptr;
logic MOSI;

endinterface
